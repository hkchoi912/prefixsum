module SparsePrefixSum(
  input          clock,
  input          reset,
  input  [15:0]  io_in,
  output [111:0] io_out
);
  assign io_out = 112'h0;
endmodule
