module SparsePrefixSum(
  input          clock,
  input          reset,
  input  [31:0]  io_in,
  output [223:0] io_out
);
  assign io_out = 224'h0;
endmodule
